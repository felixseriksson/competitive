BZh91AY&SY3|iz  �ߔPx����߰?���  P8�7�ۮv�	E2�D�ڞi'�zi2h  �4����4�SF��h 2  ��	$D<I��4 �CFF�9�14L�2da0M4����%��Q�L�4C�2� � �OX�*
�B�����ʴ6 ���
,Ķ�V�Z��,ˠ8�I/Yi6S�:_-R��9)˫Slނ���.8A�d�Qg���U O�P<��+�l�0w.��ІR7A��-�3��V���X����f�@K� 5C�f�+�6t�L�Ucd�U�k�[��a���l��<&�i_�q��¡I�����M��Tf�6r�25c�,ްF���.̻3z#Kݜ{�&�$�;�/,5�<٥�G
�Nڤ��+�>�+`榭,��
!#����GE��8}�>P�5"0�/ػ�?��
{ũ��.��B��+?,��\����{��گ�U��Ʈy/KQ��/��a~=
�٢Izy���2���	���ӮX���ELįC� ׊��d�`��\�.�M� ��,��(�v"�T,�tP[ԤI�12���
0]hrp)	Ċ�x��P �V�"XU�q���#� �tDoM�*���)��U�3�\v�Ċ�Dt��)^���!eF��7el�v���(s��)^�Zf��mn�*�ʋ �MD�K7��;�j� ͔j��Y�~4J��]�0�P�-sQ^(�@��LzF�Z*�n���a���%�HL���1���cE[�q!]x:&��^�.�q>�^��RK��F�К�<cg¡�D��>�g��h�h��khI�!<s�[�(�P�"�IeҰU����rE8P�3|iz